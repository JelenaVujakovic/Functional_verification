//------------------------------------------------------------------------------
// Copyright (c) 2020 Elsys Eastern Europe
// All rights reserved.
//------------------------------------------------------------------------------
// File name  : axi_lite_common.sv
// Developer  : Jelena Vujakovic
// Date       : Aug 8, 2020
// Description: 
// Notes      : 
//
//------------------------------------------------------------------------------

`ifndef AXI_LITE_COMMON_SV
`define AXI_LITE_COMMON_SV

typedef enum bit {
  AXI_LITE_LOW_E  = 0,
  AXI_LITE_HIGH_E = 1
} axi_lite_signal_value_e;

`endif // AXI_LITE_COMMON_SV
