`ifndef AXI_LITE_COMMON_SV
`define AXI_LITE_COMMON_SV

parameter int BLOCK_SIZE = 32768;

parameter int RESET_REG_ADDR = 0;
parameter int START_REG_ADDR = 4;
parameter int READY_REG_ADDR = 8;

`endif // AXI_LITE_COMMON_SV
