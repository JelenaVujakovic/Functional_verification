`ifndef AXI_LITE_SEQ_LIB_SV
`define AXI_LITE_SEQ_LIB_SV

`include "axi_lite_basic_seq.sv"
`include "axi_lite_write_seq.sv"
`include "axi_lite_read_seq.sv"
`include "axi_lite_read_and_write_seq.sv"

`endif // AXI_LITE_SEQ_LIB_SV
