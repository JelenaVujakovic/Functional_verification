`ifndef SCRAMBLER_IP_VIR_SEQUENCE_SV
`define SCRAMBLER_IP_VIR_SEQUENCE_SV

class scrambler_ip_vir_sequence extends scrambler_ip_base_vir;
  
	`uvm_object_utils (scrambler_ip_vir_sequence)


endclass

`endif 
