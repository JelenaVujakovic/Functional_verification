//------------------------------------------------------------------------------
// Copyright (c) 2020 Elsys Eastern Europe
// All rights reserved.
//------------------------------------------------------------------------------
// File name  : bram_a_common.sv
// Developer  : Jelena Vujakovic
// Date       : Aug 8, 2020
// Description: 
// Notes      : 
//
//------------------------------------------------------------------------------

`ifndef BRAM_A_COMMON_SV
`define BRAM_A_COMMON_SV

typedef enum bit {
  BRAM_A_LOW_E  = 0,
  BRAM_A_HIGH_E = 1
} bram_a_signal_value_e;

`endif // BRAM_A_COMMON_SV
