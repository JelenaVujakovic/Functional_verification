`ifndef BRAM_B_COMMON_SV
`define BRAM_B_COMMON_SV

parameter int BLOCK_SIZE = 8192;


`endif // BRAM_B_COMMON_SV
