//------------------------------------------------------------------------------
// Copyright (c) 2020 Elsys Eastern Europe
// All rights reserved.
//------------------------------------------------------------------------------
// File name  : bram_b_seq_lib.sv
// Developer  : Jelena Vujakovic
// Date       : Aug 8, 2020
// Description: 
// Notes      : 
//
//------------------------------------------------------------------------------

`ifndef BRAM_B_SEQ_LIB_SV
`define BRAM_B_SEQ_LIB_SV

`include "bram_b_basic_seq.sv"

`endif // BRAM_B_SEQ_LIB_SV
